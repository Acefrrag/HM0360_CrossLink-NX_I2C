library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity HM0360_Interface_tb is

end HM0360_Interface_tb;

Architecture Behavioral of HM0360_Interface_tb is

begin

end Behavioral;
