component PLL_sync_clk is
    port(
        clki_i: in std_logic;
        clkop_o: out std_logic
    );
end component;

__: PLL_sync_clk port map(
    clki_i=>,
    clkop_o=>
);
